import Ethernet::*;
import StructDefines::*;
typedef union tagged {
    struct {
    } ReqT;
    struct {
    } ReqT;
    struct {
    } ReqT;
} ForwardTblParam deriving (Bits, Eq, FShow);
import Ethernet::*;
import StructDefines::*;
