method Action forward_tbl_add_entry(ForwardTblReqT key, ForwardTblRspT val);
