
typedef enum {IfcNamesNone=0,
PlatformIfcNames_MemServerRequestS2H=1,
PlatformIfcNames_MMURequestS2H=2,
PlatformIfcNames_MemServerIndicationH2S=3,
PlatformIfcNames_MMUIndicationH2S=4,
IfcNames_MainIndicationH2S=5,
IfcNames_MemServerIndicationH2S=6,
IfcNames_MainRequestS2H=7
} IfcNames deriving (Eq,Bits);
