method forward_tbl_add_entry = prog.forward_tbl_add_entry;
